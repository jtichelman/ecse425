--Computer Org. and Arch. Project Part 2
--Tai Hung (Henry) Lu, Saki Kajita, Jeffrey Tichelman, Francois Parent
--Description: Memory controller for interacting with main memory

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

entity mem_controller is
	Generic (
		Mem_Size_in_Word : integer:=1024;	
		Num_Bytes_in_Word: integer:=4;
		Num_Bits_in_Byte: integer := 8; 
		Read_Delay: integer:=0; 
		Write_Delay:integer:=0
	);
	
	Port(
		clock : in std_logic;
		
		--Ports from IF stage
		address_if : in integer;
		read_en_if : in std_logic;
		rd_ready_if : out std_logic;
		data_if : inout std_logic_vector((Num_Bytes_in_Word*Num_Bits_in_Byte)-1 downto 0);  
		
		--Ports from MEM stage
		address_mem : in integer;
		wordbyte_mem : in std_logic;
		write_en_mem : in std_logic;
		read_en_mem : in std_logic;
		wr_done_mem : out std_logic;
		rd_ready_mem : out std_logic;
		data_mem : inout std_logic_vector((Num_Bytes_in_Word*Num_Bits_in_Byte)-1 downto 0); 
	
		--Ports to main memory
		address_out : out integer;
		word_byte_out : out std_logic;
		write_en_out : out std_logic;
		wr_done_in : in std_logic;
		read_en_out : out std_logic;
		rd_ready_in : in std_logic;
		data_inout : inout std_logic_vector((Num_Bytes_in_Word*Num_Bits_in_Byte)-1 downto 0)
	);
End mem_controller;

Architecture implementation of mem_controller is
	
	--State declarations
	type mem_state is (INPUT_STATE, READ_STATE, WRITE_STATE);
	signal current_state : mem_state := INPUT_STATE;
	
	Begin
	
	mem_process : process(clock)
	Begin
		if (clock = '1') then
			case current_state is
				--Waiting for input from either IF stage or MEM stage
				when INPUT_STATE =>
					data_if <= "ZZZZZZZZZZZZZZZZZZZZZZ";
					data_mem <= "ZZZZZZZZZZZZZZZZZZZZZZ";
					if read_en_if = '1' then	--IF read
						read_en_out <= '1';
						write_en_out <= '0';
						address_out <= address_if;
						word_byte_out <= '1';
						current_state <= READ_STATE; 
					elsif read_en_mem = '1' then		--MEM read
						read_en_out <='1';
						write_en_out <= '0';
						address_out <= address_mem;
						word_byte_out <= wordbyte_mem;
						current_state <= READ_STATE;
					elsif write_en_mem = '1' then		--MEM write
						read_en_out <='0';
						write_en_out <= '1';
						address_out <= address_mem;
						word_byte_out <= wordbyte_mem;
						current_state <= WRITE_STATE;
					else								--No memory operation
						read_en_out <='0';
						write_en_out <= '0';
						address_out <= address_mem;
						word_byte_out <= wordbyte_mem;
						current_state <= INPUT_STATE;
						data_inout <= "ZZZZZZZZZZZZZZZZZZZZZZ";
					end if;
				
				--Perform read operation on main memory
				when READ_STATE =>
					wr_done_mem<= '0';
					rd_ready_if <='0';
					rd_ready_mem <= '0';
					if (rd_ready_in = '1') then
						read_en_out <= '0';
						if (read_en_if = '1') then	-- Read to fetch
							data_if <= data_inout;
							data_mem <= "ZZZZZZZZZZZZZZZZZZZZZZ";
							rd_ready_if <= '1';
						end if;
						if (read_en_mem = '1') then	--Read to MEM
							data_mem <= data_inout;
							data_if <= "ZZZZZZZZZZZZZZZZZZZZZZ";
							rd_ready_mem <='1';
						end if;
						current_state <= INPUT_STATE;
					else 
						current_state <= READ_STATE;
					end if;
					
				--Perform write operation on main memory
				when WRITE_STATE =>
					rd_ready_if <= '0';
					rd_ready_mem <= '0';
					if (wr_done_in = '1') then
						write_en_out <= '0';
						wr_done_mem <= '1';
						current_state <= INPUT_STATE;
					else 
						current_state <= WRITE_STATE;
					end if;
				
			end case;
		end if;
	End process;

End implementation;